CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1360 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1360 728
177209362 0
0
6 Title:
5 Name:
0
0
0
26
14 Logic Display~
6 1104 297 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
0
0
8 2-In OR~
219 964 315 0 1 22
0 0
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1302252036
65 0 0 0 4 1 7 0
1 U
4441 0 0
0
0
8 4-In OR~
219 804 222 0 1 22
0 0
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0
65 0 0 0 2 2 6 0
1 U
3618 0 0
0
0
8 4-In OR~
219 807 419 0 1 22
0 0
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 1251920387
65 0 0 0 2 1 6 0
1 U
6153 0 0
0
0
13 Logic Switch~
5 383 32 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 312 32 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 242 35 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 94 529 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 95 473 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 92 415 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 91 363 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 91 294 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 94 242 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 94 185 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 96 127 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
9 Inverter~
13 420 83 0 2 22
0 4 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 5 0
1 U
4718 0 0
0
0
9 Inverter~
13 345 84 0 2 22
0 3 6
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 5 0
1 U
3874 0 0
0
0
9 Inverter~
13 266 79 0 2 22
0 2 7
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 5 0
1 U
6671 0 0
0
0
9 4-In AND~
219 616 159 0 5 22
0 14 5 6 7 16
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 2 4 0
1 U
3789 0 0
0
0
9 4-In AND~
219 617 205 0 5 22
0 15 4 6 7 17
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 1 4 0
1 U
4871 0 0
0
0
9 4-In AND~
219 616 254 0 5 22
0 13 5 3 7 18
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 2 3 0
1 U
3750 0 0
0
0
9 4-In AND~
219 616 303 0 5 22
0 12 4 3 7 19
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 1 3 0
1 U
8778 0 0
0
0
9 4-In AND~
219 616 357 0 5 22
0 11 5 6 2 20
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 2 2 0
1 U
538 0 0
0
0
9 4-In AND~
219 616 405 0 5 22
0 10 4 6 2 21
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 1 2 0
1 U
6843 0 0
0
0
9 4-In AND~
219 617 449 0 5 22
0 9 5 3 2 22
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 2 1 0
1 U
3136 0 0
0
0
9 4-In AND~
219 616 496 0 5 22
0 8 4 3 2 23
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 512 2 1 1 0
1 U
5950 0 0
0
0
51
1 3 0 0 0 0 0 1 2 0 0 5
1104 315
1104 319
1005 319
1005 315
997 315
5 2 0 0 0 0 0 4 2 0 0 4
840 419
943 419
943 324
951 324
5 1 0 0 0 0 0 3 2 0 0 4
837 222
943 222
943 306
951 306
5 3 0 0 0 0 0 26 4 0 0 4
637 496
782 496
782 424
790 424
5 3 0 0 0 0 0 25 4 0 0 4
638 449
782 449
782 424
790 424
5 2 0 0 0 0 0 24 4 0 0 4
637 405
782 405
782 415
790 415
5 1 0 0 0 0 0 23 4 0 0 4
637 357
782 357
782 406
790 406
5 3 0 0 0 0 0 22 3 0 0 4
637 303
779 303
779 227
787 227
5 3 0 0 0 0 0 21 3 0 0 4
637 254
779 254
779 227
787 227
5 2 0 0 0 0 0 20 3 0 0 4
638 205
779 205
779 218
787 218
5 1 0 0 0 0 0 19 3 0 0 4
637 159
779 159
779 209
787 209
4 0 2 0 0 4096 0 26 0 0 48 2
592 510
242 510
0 3 3 0 0 4096 0 0 26 47 0 2
312 501
592 501
2 0 4 0 0 4096 0 26 0 0 46 2
592 492
383 492
4 0 2 0 0 4096 0 25 0 0 48 2
593 463
242 463
3 0 3 0 0 16 0 25 0 0 47 3
593 454
593 455
312 455
2 0 5 0 0 4096 0 25 0 0 36 4
593 445
428 445
428 446
423 446
4 0 2 0 0 0 0 24 0 0 48 4
592 419
247 419
247 420
242 420
3 2 6 0 0 4096 0 24 17 0 0 3
592 410
348 410
348 102
2 0 4 0 0 0 0 24 0 0 46 2
592 401
383 401
4 0 2 0 0 0 0 23 0 0 48 2
592 371
242 371
3 0 6 0 0 0 0 23 0 0 19 4
592 362
588 362
588 378
348 378
2 0 5 0 0 4096 0 23 0 0 36 2
592 353
423 353
4 0 7 0 0 4096 0 22 0 0 37 4
592 317
274 317
274 318
269 318
3 0 3 0 0 0 0 22 0 0 47 4
592 308
317 308
317 309
312 309
2 0 4 0 0 0 0 22 0 0 46 2
592 299
383 299
4 0 7 0 0 4096 0 21 0 0 37 2
592 268
269 268
3 0 3 0 0 0 0 21 0 0 47 2
592 259
312 259
2 0 5 0 0 0 0 21 0 0 36 2
592 250
423 250
4 0 7 0 0 0 0 20 0 0 37 4
593 219
274 219
274 220
269 220
3 0 6 0 0 0 0 20 0 0 19 4
593 210
353 210
353 211
348 211
2 0 4 0 0 4096 0 20 0 0 46 2
593 201
383 201
4 0 7 0 0 0 0 19 0 0 37 2
592 173
269 173
0 3 6 0 0 0 0 0 19 19 0 2
348 164
592 164
2 0 5 0 0 0 0 19 0 0 36 4
592 155
428 155
428 156
423 156
2 0 5 0 0 4224 0 16 0 0 0 2
423 101
423 446
2 0 7 0 0 4224 0 18 0 0 0 2
269 97
269 318
1 1 8 0 0 4224 0 8 26 0 0 4
106 529
584 529
584 483
592 483
1 1 9 0 0 4224 0 9 25 0 0 4
107 473
585 473
585 436
593 436
1 1 10 0 0 4224 0 10 24 0 0 4
104 415
584 415
584 392
592 392
1 1 11 0 0 4224 0 11 23 0 0 4
103 363
584 363
584 344
592 344
1 1 12 0 0 4224 0 12 22 0 0 4
103 294
584 294
584 290
592 290
1 1 13 0 0 4224 0 13 21 0 0 4
106 242
584 242
584 241
592 241
1 1 14 0 0 4224 0 15 19 0 0 4
108 127
584 127
584 146
592 146
1 1 15 0 0 4224 0 14 20 0 0 4
106 185
585 185
585 192
593 192
0 0 4 0 0 4224 0 0 0 49 0 2
383 56
383 492
0 0 3 0 0 4224 0 0 0 50 0 2
312 58
312 501
0 0 2 0 0 4224 0 0 0 51 0 2
242 53
242 511
1 1 4 0 0 0 0 5 16 0 0 4
383 44
383 57
423 57
423 65
1 1 3 0 0 0 0 6 17 0 0 4
312 44
312 58
348 58
348 66
1 1 2 0 0 0 0 7 18 0 0 4
242 47
242 53
269 53
269 61
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
