CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 100 9
0 71 1359 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1359 728
177209362 0
0
6 Title:
5 Name:
0
0
0
39
13 Logic Switch~
5 491 25 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 154 30 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 317 27 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
7 Ground~
168 1303 81 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
9 3-In AND~
219 932 935 0 4 22
0 12 5 11 10
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 10 0
1 U
5394 0 0
0
0
8 4-In OR~
219 1119 800 0 5 22
0 7 8 9 10 6
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 1302252036
65 0 0 0 2 1 11 0
1 U
7734 0 0
0
0
8 3-In OR~
219 1066 286 0 4 22
0 19 18 17 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U9B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 9 0
1 U
9914 0 0
0
0
9 Inverter~
13 783 200 0 2 22
0 12 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 6 0
1 U
3747 0 0
0
0
9 3-In AND~
219 933 376 0 4 22
0 20 5 22 17
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 10 0
1 U
3549 0 0
0
0
9 CC 7-Seg~
183 1259 168 0 17 19
10 27 16 26 6 25 24 23 40 2
0 0 0 0 1 0 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
7931 0 0
0
0
8 3-In OR~
219 1092 1602 0 4 22
0 12 29 28 23
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U9A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 9 0
1 U
9325 0 0
0
0
9 2-In AND~
219 937 1577 0 3 22
0 31 13 29
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 5 0
1 U
8903 0 0
0
0
9 2-In AND~
219 936 1651 0 3 22
0 5 30 28
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 5 0
1 U
3834 0 0
0
0
8 3-In OR~
219 1092 1354 0 4 22
0 4 3 32 24
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 8 0
1 U
3363 0 0
0
0
8 3-In OR~
219 1086 1089 0 4 22
0 35 5 33 25
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 8 0
1 U
7668 0 0
0
0
8 2-In OR~
219 1087 535 0 3 22
0 38 37 26
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 7 0
1 U
4718 0 0
0
0
9 Inverter~
13 797 1661 0 2 22
0 13 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 6 0
1 U
3874 0 0
0
0
9 Inverter~
13 798 1611 0 2 22
0 5 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 6 0
1 U
6671 0 0
0
0
9 Inverter~
13 803 1456 0 2 22
0 13 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 6 0
1 U
3789 0 0
0
0
9 Inverter~
13 804 1378 0 2 22
0 5 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 6 0
1 U
4871 0 0
0
0
9 Inverter~
13 807 1308 0 2 22
0 12 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 6 0
1 U
3750 0 0
0
0
9 2-In AND~
219 935 1144 0 3 22
0 34 36 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 5 0
1 U
8778 0 0
0
0
9 Inverter~
13 804 1173 0 2 22
0 13 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 4 0
1 U
538 0 0
0
0
9 Inverter~
13 805 1098 0 2 22
0 5 34
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 4 0
1 U
6843 0 0
0
0
9 Inverter~
13 802 1023 0 2 22
0 12 35
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 4 0
1 U
3136 0 0
0
0
9 2-In AND~
219 933 853 0 3 22
0 14 13 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
5950 0 0
0
0
9 2-In AND~
219 933 778 0 3 22
0 15 13 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
5670 0 0
0
0
9 2-In AND~
219 928 704 0 3 22
0 15 14 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
6828 0 0
0
0
9 Inverter~
13 798 856 0 2 22
0 13 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 4 0
1 U
6735 0 0
0
0
9 Inverter~
13 798 788 0 2 22
0 5 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
8365 0 0
0
0
9 Inverter~
13 797 712 0 2 22
0 12 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
4132 0 0
0
0
9 Inverter~
13 783 261 0 2 22
0 5 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 6 1 0
1 U
4551 0 0
0
0
9 Inverter~
13 785 341 0 2 22
0 13 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 1 0
1 U
3635 0 0
0
0
9 2-In AND~
219 935 299 0 3 22
0 21 41 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 512 4 2 3 0
1 U
3973 0 0
0
0
9 2-In AND~
219 934 210 0 3 22
0 12 21 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
3851 0 0
0
0
9 2-In AND~
219 923 572 0 3 22
0 39 13 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 2 0
1 U
8383 0 0
0
0
9 2-In AND~
219 925 495 0 3 22
0 12 39 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 2 0
1 U
9334 0 0
0
0
9 Inverter~
13 796 526 0 2 22
0 5 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 1 0
1 U
7471 0 0
0
0
9 Inverter~
13 775 90 0 2 22
0 13 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
3334 0 0
0
0
68
2 2 3 0 0 12416 0 20 14 0 0 4
825 1378
952 1378
952 1354
1080 1354
2 1 4 0 0 4224 0 21 14 0 0 4
828 1308
1055 1308
1055 1345
1079 1345
9 1 2 0 0 4224 0 10 4 0 0 3
1259 126
1259 75
1303 75
0 2 5 0 0 8192 0 0 9 5 0 5
716 261
716 299
824 299
824 376
909 376
1 0 5 0 0 4096 0 32 0 0 66 2
768 261
317 261
5 4 6 0 0 8320 0 6 10 0 0 3
1152 800
1256 800
1256 204
3 1 7 0 0 4224 0 28 6 0 0 3
949 704
1102 704
1102 787
3 2 8 0 0 4224 0 27 6 0 0 4
954 778
1087 778
1087 796
1102 796
3 3 9 0 0 4224 0 26 6 0 0 4
954 853
1086 853
1086 805
1102 805
4 4 10 0 0 4224 0 5 6 0 0 3
953 935
1102 935
1102 814
2 3 11 0 0 8320 0 29 5 0 0 4
819 856
870 856
870 944
908 944
0 2 5 0 0 0 0 0 5 59 0 3
729 788
729 935
908 935
0 1 12 0 0 8192 0 0 5 60 0 3
693 712
693 926
908 926
0 2 13 0 0 4096 0 0 26 16 0 3
896 817
896 862
909 862
0 1 14 0 0 4096 0 0 26 18 0 3
886 788
886 844
909 844
0 2 13 0 0 8192 0 0 27 58 0 5
750 856
750 817
897 817
897 787
909 787
0 1 15 0 0 4224 0 0 27 19 0 3
869 712
869 769
909 769
2 2 14 0 0 8320 0 30 28 0 0 4
819 788
886 788
886 713
904 713
2 1 15 0 0 0 0 31 28 0 0 4
818 712
870 712
870 695
904 695
4 2 16 0 0 4224 0 7 10 0 0 3
1099 286
1244 286
1244 204
4 3 17 0 0 4224 0 9 7 0 0 4
954 376
1037 376
1037 295
1053 295
3 2 18 0 0 4224 0 34 7 0 0 4
956 299
1015 299
1015 286
1054 286
3 1 19 0 0 8320 0 35 7 0 0 4
955 210
1015 210
1015 277
1053 277
2 1 20 0 0 8320 0 8 9 0 0 4
804 200
843 200
843 367
909 367
0 1 13 0 0 8192 0 0 33 65 0 3
491 339
491 341
770 341
0 1 21 0 0 8192 0 0 34 28 0 3
879 261
879 290
911 290
0 1 12 0 0 0 0 0 35 30 0 5
716 200
716 167
880 167
880 201
910 201
2 2 21 0 0 4224 0 32 35 0 0 4
804 261
880 261
880 219
910 219
2 3 22 0 0 8320 0 33 9 0 0 3
806 341
806 385
909 385
1 0 12 0 0 4096 0 8 0 0 67 2
768 200
154 200
0 2 5 0 0 0 0 0 15 56 0 5
687 1098
687 1060
972 1060
972 1089
1074 1089
7 4 23 0 0 4224 0 10 11 0 0 3
1274 204
1274 1602
1125 1602
6 4 24 0 0 4224 0 10 14 0 0 3
1268 204
1268 1354
1125 1354
5 4 25 0 0 4224 0 10 15 0 0 3
1262 204
1262 1089
1119 1089
3 3 26 0 0 8320 0 16 10 0 0 3
1120 535
1250 535
1250 204
2 1 27 0 0 4224 0 39 10 0 0 5
796 90
1180 90
1180 218
1238 218
1238 204
3 3 28 0 0 4224 0 13 11 0 0 4
957 1651
1057 1651
1057 1611
1079 1611
3 2 29 0 0 4224 0 12 11 0 0 4
958 1577
1036 1577
1036 1602
1080 1602
0 2 13 0 0 0 0 0 12 42 0 3
698 1661
698 1586
913 1586
2 2 30 0 0 8320 0 17 13 0 0 3
818 1661
818 1660
912 1660
0 1 5 0 0 0 0 0 13 43 0 5
739 1611
739 1636
902 1636
902 1642
912 1642
0 1 13 0 0 8192 0 0 17 47 0 3
491 1456
491 1661
782 1661
0 1 5 0 0 8192 0 0 18 48 0 3
317 1378
317 1611
783 1611
2 1 31 0 0 4224 0 18 12 0 0 4
819 1611
873 1611
873 1568
913 1568
0 1 12 0 0 8320 0 0 11 49 0 5
154 1307
154 1527
1057 1527
1057 1593
1079 1593
2 3 32 0 0 4224 0 19 14 0 0 4
824 1456
1055 1456
1055 1363
1079 1363
0 1 13 0 0 8192 0 0 19 55 0 3
491 1173
491 1456
788 1456
0 1 5 0 0 8192 0 0 20 56 0 3
317 1097
317 1378
789 1378
0 1 12 0 0 0 0 0 21 57 0 3
154 1023
154 1308
792 1308
3 3 33 0 0 4224 0 22 15 0 0 6
956 1144
1032 1144
1032 1112
1062 1112
1062 1098
1073 1098
0 0 34 0 0 4224 0 0 0 53 0 2
903 1098
904 1098
2 1 35 0 0 4224 0 25 15 0 0 4
823 1023
1032 1023
1032 1080
1073 1080
2 1 34 0 0 4224 0 24 22 0 0 4
826 1098
903 1098
903 1135
911 1135
2 2 36 0 0 4224 0 23 22 0 0 4
825 1173
903 1173
903 1153
911 1153
0 1 13 0 0 4096 0 0 23 58 0 3
491 855
491 1173
789 1173
0 1 5 0 0 8320 0 0 24 59 0 3
317 786
317 1098
790 1098
0 1 12 0 0 0 0 0 25 60 0 3
154 711
154 1023
787 1023
0 1 13 0 0 0 0 0 29 65 0 3
491 579
491 856
783 856
0 1 5 0 0 0 0 0 30 66 0 3
317 526
317 788
783 788
0 1 12 0 0 0 0 0 31 67 0 3
154 486
154 712
782 712
3 2 37 0 0 4224 0 36 16 0 0 4
944 572
1032 572
1032 544
1074 544
3 1 38 0 0 4224 0 37 16 0 0 4
946 495
1031 495
1031 526
1074 526
0 1 39 0 0 4096 0 0 36 64 0 3
888 526
888 563
899 563
2 2 39 0 0 4224 0 38 37 0 0 4
817 526
888 526
888 504
901 504
0 2 13 0 0 4224 0 0 36 68 0 3
491 88
491 581
899 581
1 1 5 0 0 4224 0 3 38 0 0 3
317 39
317 526
781 526
1 1 12 0 0 0 0 2 37 0 0 3
154 42
154 486
901 486
1 1 13 0 0 0 0 1 39 0 0 3
491 37
491 90
760 90
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
